*COMPARATOR 

.param p_wp = 2.56

.SUBCKT COMP VCMP_OUT VSTORE VRAMP VBN1 VDD VSS


* Current mirror
M5 VMIRROR VMIRROR VDD VDD pmos  W = {0.65u*p_wp} L=0.13u

M6 VDM2 VMIRROR VDD VDD pmos  W = {0.65u*p_wp} L=0.13u

* Comparing VRAMP to VSTORE
M3 VMIRROR VSTORE VDM1 VSS nmos W=0.65u L=0.13u

M4 VDM2 VRAMP VDM1 VSS nmos W=0.65u L=0.13u


M1 VDM1 VBN1 VSS VSS nmos W=0.65u L=0.13u
M2 VINV VBN1 VSS VSS nmos W=0.65u L=0.13u

M7 VINV VDM2 VDD VDD pmos  W = {0.65u*p_wp} L=0.13u

*inverter
M8 VCMP_OUT VINV VDD VDD pmos W = {0.65u*p_wp} L=0.13u
M9 VCMP_OUT VINV VSS VSS nmos W=0.65u L=0.13u

.ENDS
