*MEMORY CELL

.SUBCKT MEMCELL READ VCMP_OUT IO VSS
M12 VG VCMP_OUT IO VSS nmos  w=0.2u  l=0.13u
M13 IO READ DMEM VSS nmos  w=0.4u  l=0.13u
M14 DMEM VG VSS VSS nmos  w=1u  l=0.13u
C2 VG VSS 1p
.ENDS


