*MEMORY CELL

.SUBCKT MEMCELL READ WRITE IO VSS
M1 VG WRITE IO VSS nmos  w=0.2u  l=0.13u
M2 IO READ DMEM VSS nmos  w=0.4u  l=0.13u
M3 DMEM VG VSS VSS nmos  w=0.2u  l=0.13u
C1 VG VSS 1p

.ENDS


