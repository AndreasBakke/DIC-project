*8 BITS OF MEMORY

.include memcell.cir

.SUBCKT MEMORY READ VCMP_OUT
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

XM1 READ VCMP_OUT DATA_0 VSS MEMCELL
XM2 READ VCMP_OUT DATA_1 VSS MEMCELL
XM3 READ VCMP_OUT DATA_2 VSS MEMCELL
XM4 READ VCMP_OUT DATA_3 VSS MEMCELL
XM5 READ VCMP_OUT DATA_4 VSS MEMCELL
XM6 READ VCMP_OUT DATA_5 VSS MEMCELL
XM7 READ VCMP_OUT DATA_6 VSS MEMCELL
XM8 READ VCMP_OUT DATA_7 VSS MEMCELL

.ENDS
